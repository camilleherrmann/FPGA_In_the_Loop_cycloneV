library ieee;
use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
use ieee.std_Logic_unsigned.all;

entity in_conv is 
generic(	
		NUM_CHANNEL 		: integer 	:= 40;
		CHANNEL_WIDTH		: integer 	:= 6  
	);
	port (
			clk_b    						: IN  std_logic;
			enb    							: IN  std_logic;
			reset  							: IN  std_logic;
			
			-- from SRAM B
			address_b						: OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
			data_b							: OUT STD_LOGIC_VECTOR (39 DOWNTO 0):= (others => '0');
			rden_b							: OUT STD_LOGIC  := '1';
			wren_b							: OUT STD_LOGIC  := '0';
			q_b								: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
			
			--from AST interface  
			ast_source_ready				: in std_logic; 
			ast_source_channel			: in std_logic_vector(CHANNEL_WIDTH-1 downto 0);
	
			--to AST interface
			ast_sink_valid					: out std_logic;													 												
			ast_sink_sop					: out std_logic;													 
			ast_sink_eop					: out std_logic;	
			ast_sink_ready					: out std_logic; 
			ast_sink_data					: out std_logic_vector(31 downto 0);
			ast_sink_channel				: out std_logic_vector(CHANNEL_WIDTH-1 downto 0)	
		);
end entity in_conv;

architecture behav of in_conv is

type 	 states								is (state1, state2);
signal state								: states;
signal s_channel 							: std_logic_vector(CHANNEL_WIDTH-1 downto 0);
signal s_sop, s_eop,s_valid, s_rden : std_logic;
signal addr 								: std_logic_vector(9 downto 0);
signal out_ready 							: std_logic;
signal round1								: std_logic_vector(1 downto 0):="00";
signal round2 								: std_logic_vector(7 downto 0):=(others => '0');

begin

	u_readenable : process(reset,enb)
	begin
		if (reset = '0') then
			s_rden	  				<='0';		
			elsif (enb = '1')  then
				s_rden				<='1';
		end if;
	end process;
	
	u_ast_valid : process (clk_b,reset,enb)
		begin
			if (reset = '0') then
			s_valid 					<= '0';		
			elsif(clk_b'event and clk_b='1') then
				if (s_rden = '1') then 
					s_valid 			<='1';
				else 	s_valid		<= '0';
				end if;
			end if;
	end process;
			


	u_main_part : process(reset,clk_b)
	begin
		if (reset = '0') then
			state 				<= state1;
			s_channel			<= (others => '0');
			out_ready			<= '0';
			s_sop 				<= '0';
			s_eop					<= '0';
		
		elsif (clk_b'event and clk_b='1') then
		
		case state is 
		
			when state1 =>
				out_ready 		<= '1';
				s_eop				<= '0';
				if (s_valid = '1' and ast_source_ready = '1') then
				   out_ready	<= '0';
					s_sop			<= '1';
					s_channel 	<= ast_source_channel;
					state			<= state2;
				end if;
			
			when state2 =>
				s_sop 			<= '0';
				if(s_valid = '1' and ast_source_ready = '1') then 
				s_eop				<= '1';
				out_ready		<= '1';
				state				<= state1;
				end if;
				
			when others =>
				out_ready		<= '1';
				state				<= state1;
		end case;	
		end if;	
	end process;
	
	u_ast_data : process(clk_b, reset, enb)
	begin
		if (reset = '0') then
			addr	  				<= (others => '0');	
			round1					<= (others => '0');	
			elsif(clk_b'event and clk_b='1') then
				if (state = state1) then 
				ast_sink_data <= q_b(31 downto 0);
				addr 	<= round1 & round2;
				round2 <= round2 + 1;
				end if;
				if (round2 = "11111111" ) then
					round1 			<= round1 + 1;
				end if;
		end if;
	end process;
			
--			
--	u_ready : process(clk_b,reset, enb)
--	begin
--		if(reset='0')then
--			out_ready	<= '0';
--		elsif(clk_b'event and clk_b='1') then
--			if (enb = '1' and in_ready ='1') then
--				out_ready <= '1';	
--			end if;
--		end if;
--	end process;
		
--	u_ast_sop : process(clk_b, reset)
--	begin
--		if (reset = '0') then
--			s_sop 					<= '0';
--		elsif(clk_b'event and clk_b='1') then
--			if (s_channel + 1 = (s_channel'range => '0')) then
--				s_sop 				<= '1';
--			else s_sop				<= '0';
--			end if;
--		end if;
--	end process;	
--		
--	u_ast_eop : process(clk_b, reset)
--	begin
--		if (reset = '0') then
--			s_eop 					<= '0';
--		elsif(clk_b'event and clk_b='1') then
--			if (s_channel + 1 = (s_channel'range => '1')) then
--				s_eop 				<= '1';
--			else s_eop				<= '0';
--			end if;
--		end if;
--	end process;
--	
--	
--	u_channel : process(clk_b, reset)
--	begin
--		if (reset = '0') then
--			s_channel 				<= (others => '0');
--		elsif (clk_b'event and clk_b='1') then
--			if (out_ready ='1' and s_valid ='1' and s_channel /= ast_source_channek) then 
--			s_channel				<= s_channel + 1;
--			end if;
--		end if;
--	end process;



	


ast_sink_channel		 <= s_channel;
ast_sink_sop			 <= s_sop;
ast_sink_eop			 <= s_eop;
ast_sink_valid			 <= s_valid;
rden_b 					 <= s_rden;
address_b 				 <= addr;
ast_sink_ready 		 <= out_ready;
	
end behav;		
			
			
			
			
			
			